package config;
    parameter ERR_STATUS_ADDRESS = 1;
    parameter PAYLOAD_ADDRESS = 2;
    parameter DATA_SIZE_ADDRESS = 4;
endpackage;